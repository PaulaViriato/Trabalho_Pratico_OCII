module banco_registradores (
input[15:0]      entrada 1,
input[15:0]      entrada 2,
output reg[31:0] saida
);

	always@(posedge clk)
	begin

	end
	
endmodule